architecture RTL1 of c is
	
begin

end architecture RTL1;