architecture RTL1 of a is
	
begin

end architecture RTL1;