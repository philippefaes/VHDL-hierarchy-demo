library ieee;
use ieee.std_logic_1164.all;

entity a is
	port (
		x : in std_logic;
		y : out std_logic
	);
end entity a;
