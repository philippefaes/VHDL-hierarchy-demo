architecture RTL2 of c is
	
begin

end architecture RTL2;
