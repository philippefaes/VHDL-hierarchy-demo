library ieee;
use ieee.std_logic_1164.all;

entity a is
	port (
		x : in std_logic;
		y : out std_logic
	);
end entity a;

architecture RTL1 of a is
	
begin

end architecture RTL1;

architecture RTL2 of a is
	
begin

end architecture RTL2;
