library ieee;
use ieee.std_logic_1164.all;

entity c is
	port (
		x : out std_logic;
		y : in std_logic
	);
end entity c;
