architecture RTL2 of a is
	
begin

end architecture RTL2;
