architecture RTL1 of b is
	
begin

end architecture RTL1;